class ptc_transaction extends uvm_sequence_item;

  rand bit [31:0] addr;
  rand bit [31:0] data; //read or write from DUT
  rand bit write; //write=1 read=0
  rand bit use_capt; // if 1 pulse the ptc_capt signal
  rand bit use_ecgt; // if set to 1, apply ptc_ecgt with value specified below
  rand bit ecgt_val; //value to be applied on ptc_ecgt (1 = high, 0 = low)

  `uvm_object_utils(ptc_transaction)

  function new(string name = "ptc_transaction");
    super.new(name);
  endfunction

  function void do_print(uvm_printer printer);
    super.do_print(printer);
    `uvm_info("PTC_TX", $sformatf(
      "\nAddress     = 0x%0h\nWrite?      = %0b\nData        = 0x%0h\nUse Capt?   = %0b\nUse ECGT?   = %0b\nECGT Value  = %0b",
      addr, write, data, use_capt, use_ecgt, ecgt_val
    ), UVM_LOW)
  endfunction

endclass